module multiply_fixed_point(
    input wire signed [15:0] integer_input,    // Số nguyên 16-bit
    input wire signed [31:0] real_input,       // Số thực 32-bit, 1 bit dấu, 3 bit nguyên, 28 bit thập phân
    output wire signed [47:0] result   // Đầu ra số nguyên 16-bit
);

// Thực hiện phép nhân, kết quả tạm thời l�  48-bit để đảm bảo không mất mát thông tin
wire signed [47:0] multiply_result = $signed(integer_input) * real_input;

// Scale v�  l� m tròn kết quả để phù hợp với đầu ra 16-bit.
// Lưu ý: Việc dịch 28 bit giúp loại bỏ phần thập phân, nhưng cần xem xét cẩn thận cách l� m tròn
//wire signed [15:0] rounded_result = multiply_result[47:28] + {{15{multiply_result[27]}}, multiply_result[27]};

assign result = multiply_result;

endmodule

`timescale 1ns / 1ps

module testbench;

    // Inputs
    reg signed [15:0] integer_input;
    reg signed [31:0] real_input;

    // Output
    wire signed [15:0] result;

    // Instantiate the Device Under Test (DUT)
    multiply_fixed_point dut (
        .integer_input(integer_input), 
        .real_input(real_input), 
        .result(result)
    );

    // Initialize all inputs
    initial begin
        // Initialize Inputs
        integer_input = 0;
        real_input = 0;

        // Wait for 100 ns for global reset to finish
        #100;
        
        // Input test values
        integer_input = 16'd17527;             // Positive integer
        real_input = 32'h007537fb;          // Positive real (1.0 in fixed-point)
        #10;                                   // Wait for the result
        
        integer_input = -16'sd1000;            // Negative integer
        real_input = -32'sd2000000000;         // Negative real (-2.0 in fixed-point)
        #10;

        integer_input = 16'sd500;             // Smaller positive integer
        real_input = 32'sd500000000;          // Smaller real (0.5 in fixed-point)
        #10;

        integer_input = -16'sd500;            // Negative integer
        real_input = 32'sd1073741824;         // Positive real approx. (0.25 in fixed-point)
        #10;
        
        integer_input = 16'sd32767;           // Max positive integer
        real_input = 32'sd1073741824;         // Real input (0.25 in fixed-point)
        #10;
        
        integer_input = -16'sd32768;          // Max negative integer
        real_input = -32'sd2147483648;        // Real input (-2.0 in fixed-point)
        #10;

        // Test rounding
        integer_input = 16'sd123;             // Test rounding
        real_input = 32'sd234881024;          // Close to 0.055 in fixed-point
        #10;

        // Complete the test
        $finish;
    end
    
    // Monitor changes and display them
    initial begin
        $monitor("At time %t, input = %d, real_input = %d, result = %d",
                 $time, integer_input, real_input, result);
    end

endmodule
