module Sign_mag_add
#(
    parameter N=4;
)