module coeffs(
	
);

endmodule