module IIR_fillter #(
	parameter DATA_BIT_NUM = 16,
	parameter DATA_BIT_NUMK = 48
)(
	input clk,
	input rst_n,
	input signed [31:0] coeff_in_1,
	input signed [31:0] coeff_in_2,
	input signed [31:0] coeff_in_3,
	input signed [31:0] coeff_out_1,
	input signed [31:0] coeff_out_2,
	input signed [DATA_BIT_NUM-1:0] data_in,
	output wire signed [DATA_BIT_NUM-1:0] data_out
);
wire signed [DATA_BIT_NUMK-1:0] delay_1_b;
wire signed [DATA_BIT_NUMK-1:0] delay_2_b;
reg signed [DATA_BIT_NUMK-1:0] delay_1_a;
reg signed [DATA_BIT_NUMK-1:0] delay_2_a;
wire signed [DATA_BIT_NUMK-1:0] data_in_coeff_1;
wire signed [DATA_BIT_NUMK-1:0] data_in_coeff_2;
wire signed [DATA_BIT_NUMK-1:0] data_in_coeff_3;
wire signed [DATA_BIT_NUMK-1:0] data_out_coeff_1;
wire signed [DATA_BIT_NUMK-1:0] data_out_coeff_2;
wire signed [DATA_BIT_NUMK-1:0] data_out_pre;
multiply_fixed_point multi(
	.integer_input(data_in),
	.real_input(coeff_in_1),
	.result(data_in_coeff_1)
);
multiply_fixed_point multi_1(
	.integer_input(data_in),
	.real_input(coeff_in_2),
	.result(data_in_coeff_2)
);
multiply_fixed_point multi_2(
	.integer_input(data_in),
	.real_input(coeff_in_3),
	.result(data_in_coeff_3)
);
multiply_fixed_point multi_3(
	.integer_input(data_out),
	.real_input(coeff_out_1),
	.result(data_out_coeff_1)
);
multiply_fixed_point multi_4(
	.integer_input(data_out),
	.real_input(coeff_out_2),
	.result(data_out_coeff_2)
);
assign delay_1_b=data_in_coeff_2-data_out_coeff_1+delay_2_a;
assign delay_2_b=data_in_coeff_3-data_out_coeff_2;
always@(posedge clk or negedge rst_n) begin
	if(~rst_n) begin
	delay_1_a<=0;
	delay_2_a<=0;
	end
	else begin
	delay_1_a<=delay_1_b;
	delay_2_a<=delay_2_b;
	end
end
assign data_out_pre=delay_1_a+data_in_coeff_1;
wire signed [15:0] data_out_pre_1 = data_out_pre[47:28] + {{15{data_out_pre[27]}}, data_out_pre[27]};
assign data_out=data_out_pre_1;
endmodule 
`timescale 1ns / 1ps

module testbench_1;

    // Parameters
    parameter DATA_BIT_NUM = 16;
    integer i;
    parameter SAMPLES = 1024;
    reg [DATA_BIT_NUM-1:0] data_array [0:SAMPLES-1];
    // Inputs
    reg clk;
    reg rst_n;
    reg signed [31:0] coeff_in_1;
    reg signed [31:0] coeff_in_2;
    reg signed [31:0] coeff_in_3;
    reg signed [31:0] coeff_out_1;
    reg signed [31:0] coeff_out_2;
    reg signed [DATA_BIT_NUM-1:0] data_in;

    // Outputs
    wire signed [DATA_BIT_NUM-1:0] data_out;

    // Instantiate the Unit Under Test (UUT)
    IIR_fillter #(
        .DATA_BIT_NUM(DATA_BIT_NUM)
    ) uut (
        .clk(clk), 
        .rst_n(rst_n), 
        .coeff_in_1(coeff_in_1), 
        .coeff_in_2(coeff_in_2), 
        .coeff_in_3(coeff_in_3), 
        .coeff_out_1(coeff_out_1), 
        .coeff_out_2(coeff_out_2), 
        .data_in(data_in), 
        .data_out(data_out)
    );

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk;  // Generate a clock with a period of 10 ns
    end

    // Initial Conditions and Stimuli
    initial begin
        // Initialize Inputs
        rst_n = 0;
        coeff_in_1 = 32'h000000bb; // 1.0 in fixed-point
        coeff_in_2 = 32'h00000176; // 0.5 in fixed-point
        coeff_in_3 = 32'h000000bb; // 0.25 in fixed-point
        coeff_out_1 = 32'he173bc58; // -0.5 in fixed-point
        coeff_out_2 = 32'h0e978a34; // -0.25 in fixed-point
        data_in = 0;

        // Reset the system
        #20;
        rst_n = 1;

    $readmemb("sin_noise.txt", data_array);
    #20 rst_n = 1;  // Reset deactivation aligned with the clock edge

    for (i = 0; i < SAMPLES; i = i + 1) begin
        @ (posedge clk);
        data_in = data_array[i];
    end

        // Complete the simulation
        $finish;
    end

    // Monitor changes and display them
    initial begin
        $monitor("At time %t, input = %d, output = %d",
                 $time, data_in, data_out);
    end

endmodule
